*AXA2

.subckt AXA2 a b cin sum cout vdd
*PMOS
    Mp1 vdd a sc1 a pmos_nvt l=len nfins=n
    Mp2 sc1 b sum b pmos_nvt l=len nfins=n
    Mp3 cin sum cout sum pmos_nvt l=len nfins=n
*NMOS
    Mn1 sum b a b nmos_nvt l=len nfins=n
    Mn2 sum a b a nmos_nvt l=len nfins=n
    Mn3 a sum cout sum nmos_nvt l=len nfins=n
.ends
