*circuit - SMA
.subckt SMA a b cin sum cout vdd gnd
*DUT
    *PMOS
        Mp1 vdd b sc1 vdd pmos_rvt l=len nfins=n
        Mp2 sc1 cin co vdd pmos_rvt l=len nfins=n
        Mp3 vdd b sc2 vdd pmos_rvt l=len nfins=n
        Mp4 sc2 a co vdd pmos_rvt l=len nfins=n
        Mp5 vdd a sc3 vdd pmos_rvt l=len nfins=n
        Mp6 vdd b sc3 vdd pmos_rvt l=len nfins=n
        Mp7 sc3 co su vdd pmos_rvt l=len nfins=n
        Mp8 vdd cin su vdd pmos_rvt l=len nfins=n
    *NMOS
        Mn1 co cin sd1 cin nmos_rvt l=len nfins=n
        Mn2 sd1 a gnd a nmos_rvt l=len nfins=n
        Mn3 co b gnd b nmos_rvt l=len nfins=n
        Mn4 su co sd2 co nmos_rvt l=len nfins=n
        Mn5 sd2 cin gnd cin nmos_rvt l=len nfins=n
        Mn6 su cin se1 cin nmos_rvt l=len nfins=n
        Mn7 se1 a se2 a nmos_rvt l=len nfins=n
        Mn8 se2 b gnd b nmos_rvt l=len nfins=n
    *inverter for output
        Xsum su sum vdd gnd Inv
        Xcout co cout vdd gnd Inv
.ends
