*AMA2 test COUT

*model
.include 7nm_FF.pm

*param
.param vdd = 0.7V
.param len = 7nm
.param n = 3
.param m = 1ns
.option post = 2
*sets format to .csv file
.option measform= 3
*outputs all measures to one file
.option measfile = 1


*sources
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd
*test sources
Va a_in gnd PWL('0*m' 0 '1*m' 0 '1.1*m' vdd '2*m' vdd '2.1*m' 0 '4*m' 0 '4.1*m' vdd '5*m' vdd '5.1*m' 0 '7*m' 0 '7.1*m' vdd '8*m' vdd '8.1*m' 0 '10*m' 0 '10.1*m' vdd '11*m' vdd '11.1*m' 0)
Vb b_in gnd PWL('0*m' 0 '6*m' 0 '6.1*m' vdd)
Vcin c_in gnd PWL('0*m' 0 '3*m' 0 '3.1*m' vdd '6*m' vdd '6.1*m' 0 '9*m' 0 '9.1*m' vdd)

.include INVERTER.cir
.include AMA2.cir

*IN fanout
Xinv1 a_in a_in1 vdd1 Inv
Xinv2 a_in1 a vdd1 Inv

Xinv3 b_in b_in1 vdd1 Inv
Xinv4 b_in1 b vdd1 Inv

Xinv5 c_in c_in1 vdd1 Inv
Xinv6 c_in1 cin vdd1 Inv

*****************DUT******************
XDUT a b cin sum cout vdut AMA2

*OUT fanout
Xinv8 sum sum_1 vdd2 Inv M=2
Xinv9 sum_1 sum_2 vdd2 Inv M=2

Xinv10 cout cout_1 vdd2 Inv M=2
Xinv11 cout_1 cout_2 vdd2 Inv M=2

*Measures atraso
.measure tran tplh_A00 trig v(A) val='0.5*vdd' rise=1 targ v(cout) val='0.5*vdd' rise=1
.measure tran tplh_A01 trig v(A) val='0.5*vdd' rise=2 targ v(cout) val='0.5*vdd' rise=2
.measure tran tplh_A10 trig v(A) val='0.5*vdd' rise=3 targ v(cout) val='0.5*vdd' rise=3
.measure tran tplh_A11 trig v(A) val='0.5*vdd' rise=4 targ v(cout) val='0.5*vdd' rise=4
.measure tran tphl_A00 trig v(A) val='0.5*vdd' fall=1 targ v(cout) val='0.5*vdd' fall=1
.measure tran tphl_A01 trig v(A) val='0.5*vdd' fall=2 targ v(cout) val='0.5*vdd' fall=2
.measure tran tphl_A10 trig v(A) val='0.5*vdd' fall=3 targ v(cout) val='0.5*vdd' fall=3
.measure tran tphl_A11 trig v(A) val='0.5*vdd' fall=4 targ v(cout) val='0.5*vdd' fall=4
*Measures energia
.measure tran e_in integ i(Vvdd1) from='0*m' to='12*m'
.measure tran e_fa integ i(Vvdut) from='0*m' to='12*m'
.measure tran e_out integ i(Vvdd2) from='0*m' to='12*m'

*simulation
.tran '0.1*m' '12*m

.end
