*AXA3 test SUM

*model
.include 7nm_FF.pm

*param
.param vdd = 0.7V
.param n = 3
.param m = 1n
.option post = 2
*sets format to .csv file
.option measform= 3
*outputs all measures to one file
.option measfile = 1

*sources
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd
*Vboost boost gnd 0.9V
*test sources
Va a_in gnd PWL('0*m' 0 '4.0*m' 0 '4.1*m' vdd '8.0*m' vdd '8.1*m' 0 '9.0*m' 0 '9.1*m' vdd '11.0*m' vdd '11.1*m' 0)
Vb b_in gnd PWL('0*m' 0 '2.0*m' 0 '2.1*m' vdd '3.0*m' vdd '3.1*m' 0 '5.0*m' 0 '5.1*m' vdd '10.0*m' vdd '10.1*m' 0)
Vcin c_in gnd PWL('0*m' 0 '1.0*m' 0 '1.1*m' vdd '6.0*m' vdd '6.1*m' 0 '7.0*m' 0 '7.1*m' vdd '12.0*m' vdd '12.1*m' 0)

.include INVERTER.cir
.include AXA3.cir

*IN
Xinv1 a_in a_in1 vdd1 Inv
*Xinv2 a_in1 a boost Inv
Xinv2 a_in1 a vdd1 Inv

Xinv3 b_in b_in1 vdd1 Inv
Xinv4 b_in1 b vdd1 Inv

Xinv5 c_in c_in1 vdd1 Inv
Xinv6 c_in1 cin vdd1 Inv

***************DUT******************
XDUT a b cin sum cout vdut AXA3

*OUT
Csum sum gnd 10f
Ccout cout gnd 10f

*delay
.measure tran tplh_00C trig v(Cin) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' rise=1
.measure tran tplh_0B1 trig v(B) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' rise=2
.measure tran tplh_1B1 trig v(B) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' rise=3
.measure tran tplh_11C trig v(Cin) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' rise=4
.measure tran tplh_A11 trig v(A) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' rise=5
.measure tran tplh_A01 trig v(A) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' rise=6
.measure tran tphl_0B1 trig v(B) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' fall=1
.measure tran tphl_A01 trig v(A) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' fall=2
.measure tran tphl_11C trig v(Cin) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' fall=3
.measure tran tphl_A11 trig v(A) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' fall=4
.measure tran tphl_1B1 trig v(B) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' fall=5
.measure tran tphl_00C trig v(Cin) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' fall=6

*energy
.measure tran e_in integ i(Vvdd1) from=0n to='13*m'
.measure tran e_fa integ i(Vvdut) from=0n to='13*m'
.measure tran e_out integ i(Vvdd2) from=0n to='13*m'
*.measure tran e_boost integ i(Vboost) from=0n to='13*m'

*simulation
.tran '0.1*m' '13*m'

.end
