*EXA test cout

*model
.include 7nm_FF.cir

*param
.param vdd = 0.7V
.param len = 7nm
.param n = 3
.param m = 1n
.option post = 2
*sets format to .csv file
.option measform= 3
*outputs all measures to one file
.option measfile = 1


*source
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd
*Vboost boost gnd 0.9V
*test source
Va a_in gnd PWL('0*m' 0 '3*m' 0 '3.1*m' vdd '6*m' vdd '6.1*m' 0 '9*m' 0 '9.1*m' vdd '12*m' vdd '12.1*m' 0)
Vb b_in gnd PWL('0*m' 0 '1*m' 0 '1.1*m' vdd '2*m' vdd '2.1*m' 0 '5*m' 0 '5.1*m' vdd '10*m' vdd '10.1*m' 0)
Vcin c_in gnd PWL('0*m' vdd '4*m' vdd '4.1*m' 0 '7*m' 0 '7.1*m' vdd '8*m' vdd '8.1*m' 0 '11*m' 0 '11.1*m' vdd)

.include INVERTER.cir
.include EXA.cir

*IN
Xinv1 a_in a_in1 vdd1 gnd Inv
*Xinv2 a_in1 a boost gnd Inv
Xinv2 a_in1 a vdd1 gnd Inv

Xinv3 b_in b_in1 vdd1 gnd Inv
Xinv4 b_in1 b vdd1 gnd Inv

Xinv5 c_in c_in1 vdd1 gnd Inv
Xinv6 c_in1 cin vdd1 gnd Inv

***************DUT******************
XDUT a b cin sum cout vdut gnd EXA

*OUT
Xinv7 sum  sum_1 vdd2 gnd Inv M=2
Xinv8 sum_1  sum_2 vdd2 gnd Inv M=2
Xinv9 cout cout_1 vdd2 gnd Inv M=2
Xinv10 cout_1 cout_2 vdd2 gnd Inv M=2


*Measures atraso
.measure tran tplh_0B1 trig v(B) val='0.5*vdd' rise=1 targ v(cout) val='0.5*vdd' rise=1
.measure tran tphl_0B1 trig v(B) val='0.5*vdd' fall=1 targ v(cout) val='0.5*vdd' fall=1
.measure tran tplh_A01 trig v(A) val='0.5*vdd' rise=1 targ v(cout) val='0.5*vdd' rise=2
.measure tran tphl_A01 trig v(A) val='0.5*vdd' fall=2 targ v(cout) val='0.5*vdd' fall=6
.measure tran tplh_01C trig v(Cin) val='0.5*vdd' rise=1 targ v(cout) val='0.5*vdd' rise=4
.measure tran tphl_01C trig v(Cin) val='0.5*vdd' fall=2 targ v(cout) val='0.5*vdd' fall=4
.measure tran tplh_A10 trig v(A) val='0.5*vdd' rise=2 targ v(cout) val='0.5*vdd' rise=5
.measure tran tphl_A10 trig v(A) val='0.5*vdd' fall=1 targ v(cout) val='0.5*vdd' fall=3
.measure tran tplh_1B0 trig v(B) val='0.5*vdd' rise=2 targ v(cout) val='0.5*vdd' rise=3
.measure tran tphl_1B0 trig v(B) val='0.5*vdd' fall=2 targ v(cout) val='0.5*vdd' fall=5
.measure tran tplh_10C trig v(Cin) val='0.5*vdd' rise=2 targ v(cout) val='0.5*vdd' rise=6
.measure tran tphl_10C trig v(Cin) val='0.5*vdd' fall=1 targ v(cout) val='0.5*vdd' fall=2

*Measures energia
.measure tran e_in integ i(Vvdd1) from=0n to='13*m'
.measure tran e_fa integ i(Vvdut) from=0n to='13*m'
.measure tran e_out integ i(Vvdd2) from=0n to='13*m'
.measure tran e_boost integ i(Vboost) from=0n to='13*m'

*Simulação transiente
.tran '0.1*m' '13*m'

.end
