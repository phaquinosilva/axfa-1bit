*MIRROR test SUM

*model
.include 7nm_FF.pm

*param
.param vdd = 0.7V
.param len = 7nm
.param n = 3
.param m = 1n
.option post = 2
*sets format to .csv file
.option measform= 3
*outputs all measures to one file
.option measfile = 1

*sources
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd
*sources sum
Va a_in gnd PWL('0*m' 0 '5*m' 0 '5.1*m' vdd '7*m' vdd '7.1*m' 0 '10*m' 0 '10.1*m' vdd '13*m' vdd '13.1*m' 0 '16*m' 0 '16.1*m' vdd '18*m' vdd '18.1*m' 0 '19*m' 0 '19.1*m' vdd '24*m' vdd '24.1*m' 0)
Vb b_in gnd PWL('0*m' 0 '3*m' 0 '3.1*m' vdd '4*m' vdd '4.1*m' 0 '8*m' 0 '8.1*m' vdd '9*m' vdd '9.1*m' 0 '12*m' 0 '12.1*m' vdd '20*m' vdd '20.1*m' 0 '21*m' 0 '21.1*m' vdd '23*m' vdd '23.1*m' 0)
Vcin c_in gnd PWL('0*m' 0 '1*m' 0 '1.1*m' vdd '2*m' vdd '2.1*m' 0 '6*m' 0 '6.1*m' vdd '11*m' vdd '11.1*m' 0 '14*m' 0 '14.1*m' vdd '15*m' vdd '15.1*m' 0 '17*m' 0 '17.1*m' vdd '22*m' vdd '22.1*m' 0)

.include INVERTER.cir
.include MIRROR.cir

*IN fanout
Xinv1 a_in a_in1 vdd1 gnd Inv
Xinv2 a_in1 a vdd1 gnd Inv

Xinv3 b_in b_in1 vdd1 gnd Inv
Xinv4 b_in1 b vdd1 gnd Inv

Xinv5 c_in c_in1 vdd1 gnd Inv
Xinv6 c_in1 cin vdd1 gnd Inv

*****************DUT******************
XDUT a b cin sum cout vdut gnd MIR

*OUT fanout
Xinv8 sum sum_1 vdd2 gnd Inv M=2
Xinv9 sum_1 sum_2 vdd2 gnd Inv M=2

Xinv10 cout cout_1 vdd2 gnd Inv M=2
Xinv11 cout_1 cout_2 vdd2 gnd Inv M=2

*Measures atraso
.measure tran tplh_00C trig v(Cin) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' rise=1
.measure tran tphl_00C trig v(Cin) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' fall=1
.measure tran tplh_0B0 trig v(B) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' rise=2
.measure tran tphl_0B0 trig v(B) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' fall=2
.measure tran tplh_A00 trig v(A) val='0.5*vdd' rise=1 targ v(sum) val='0.5*vdd' rise=3
.measure tran tphl_A00 trig v(A) val='0.5*vdd' fall=4 targ v(sum) val='0.5*vdd' fall=12
.measure tran tplh_0B1 trig v(B) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' rise=5
.measure tran tphl_0B1 trig v(B) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' fall=4
.measure tran tplh_01C trig v(Cin) val='0.5*vdd' fall=3 targ v(sum) val='0.5*vdd' rise=8
.measure tran tphl_01C trig v(Cin) val='0.5*vdd' rise=3 targ v(sum) val='0.5*vdd' fall=7
.measure tran tplh_A11 trig v(A) val='0.5*vdd' rise=4 targ v(sum) val='0.5*vdd' rise=10
.measure tran tphl_A11 trig v(A) val='0.5*vdd' fall=3 targ v(sum) val='0.5*vdd' fall=9
.measure tran tplh_A01 trig v(A) val='0.5*vdd' fall=1 targ v(sum) val='0.5*vdd' rise=4
.measure tran tphl_A01 trig v(A) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' fall=5
.measure tran tplh_10C trig v(Cin) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' rise=6
.measure tran tphl_10C trig v(Cin) val='0.5*vdd' rise=2 targ v(sum) val='0.5*vdd' fall=3
.measure tran tplh_1B1 trig v(B) val='0.5*vdd' rise=4 targ v(sum) val='0.5*vdd' rise=11
.measure tran tphl_1B1 trig v(B) val='0.5*vdd' fall=3 targ v(sum) val='0.5*vdd' fall=10
.measure tran tplh_A10 trig v(A) val='0.5*vdd' fall=2 targ v(sum) val='0.5*vdd' rise=7
.measure tran tphl_A10 trig v(A) val='0.5*vdd' rise=3 targ v(sum) val='0.5*vdd' fall=8
.measure tran tplh_1B0 trig v(B) val='0.5*vdd' fall=4 targ v(sum) val='0.5*vdd' rise=12
.measure tran tphl_1B0 trig v(B) val='0.5*vdd' rise=3 targ v(sum) val='0.5*vdd' fall=6
.measure tran tplh_11C trig v(Cin) val='0.5*vdd' rise=4 targ v(sum) val='0.5*vdd' rise=9
.measure tran tphl_11C trig v(Cin) val='0.5*vdd' fall=4 targ v(sum) val='0.5*vdd' fall=11

*Measures energia
.measure tran e_in integ i(Vvdd1) from=0n to='25*m'
.measure tran e_fa integ i(Vvdut) from=0n to='25*m'
.measure tran e_out integ i(Vvdd2) from=0n to='25*m'

*Simulação transiente
.tran '0.1*m' '25*m'

.end
