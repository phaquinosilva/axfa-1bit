*circuit - AXA2
.subckt AXA2 a b cin sum cout vdd
*PMOS
    Mp1 vdd a sc1 a pmos_rvt nfin=n
    Mp2 sc1 b sum b pmos_rvt nfin=n
    Mp3 cin sum cout sum pmos_rvt nfin=n
*NMOS
    Mn1 sum b a b nmos_rvt nfin=n
    Mn2 sum a b a nmos_rvt nfin=n
    Mn3 a sum cout sum nmos_rvt nfin=n
.ends
